*.subckt sar_logic clk rstn en comp cal valid result.0 result.1 result.2 result.3 result.4 result.5 sample ctlp.0 ctlp.1 ctlp.2 ctlp.3 ctlp.4 ctlp.5 ctln.0 ctln.1 ctln.2 ctln.3 ctln.4 ctln.5 trim.0 trim.1 trim.2 trim.3 trim.4 trimb.0 trimb.1 trimb.2 trimb.3 trimb.4 clkc
.subckt sarlogic on clk comp result.0 result.1 result.2 result.3 result.4 result.5 sample ctlp.0 ctlp.1 ctlp.2 ctlp.3 ctlp.4 ctlp.5 ctln.0 ctln.1 ctln.2 ctln.3 ctln.4 ctln.5 clkc 
X0 rstn 1 NOT
X1 en 2 NOT
X2 cal_itt.1 3 NOT
X3 cal_itt.2 4 NOT
X4 cal_itt.3 5 NOT
X5 comp 6 NOT
X6 cal_count.2 7 NOT
X7 cal_count.3 8 NOT
X8 en_co_clk 9 NOT
X9 trim_mask.0 10 NOT
X10 trim_val.4 11 NOT
X11 state.0 12 NOT
X12 state.1 13 NOT
X13 state.2 14 NOT
X14 result.0 15 NOT
X15 result.1 16 NOT
X16 result.2 17 NOT
X17 result.3 18 NOT
X18 result.4 19 NOT
X19 result.5 20 NOT
*X20 result.6 21 NOT
*X21 result.7 22 NOT
*X22 result.8 23 NOT
*X23 result.9 24 NOT
X24 state.0 state.1 25 NOR
X25 state.2 25 26 NAND
X26 26 valid NOT
X27 state.0 state.2 27 NOR
X28 27 28 NOT
X29 state.1 27 29 NAND
X30 29 30 NOT
X31 12 state.1 31 NOR
X32 state.0 13 32 NAND
X33 14 32 33 NOR
X34 state.2 31 34 NAND
X35 29 34 sample NAND
X36 cal_itt.0 cal_itt.1 35 NAND
X37 35 36 NOT
X38 4 35 37 NOR
X39 cal_itt.2 36 38 NAND
X40 cal_itt.3 38 39 NOR
X41 5 37 40 NAND
X42 10 40 41 NOR
X43 trim_mask.0 39 42 NAND
X44 cal_itt.0 42 43 NAND
X45 33 43 44 NAND
X46 en state.2 45 NOR
X47 45 46 NOT
X48 32 45 47 NOR
X49 31 46 48 NAND
X50 cal_itt.0 48 49 NAND
X51 44 49 50.0 NAND
X52 cal_itt.0 cal_itt.1 51 NOR
X53 3 47 52 NOR
X54 35 41 53 NOR
X55 34 53 54 NOR
X56 52 54 55 NOR
X57 51 55 50.1 NOR
X58 4 35 56 NAND
X59 38 56 57 NAND
X60 42 57 58 NAND
X61 33 58 59 NAND
X62 cal_itt.2 48 60 NAND
X63 59 60 50.2 NAND
X64 12 state.2 61 NOR
X65 61 62 NOT
X66 state.2 32 63 NOR
X67 63 64 NOT
X68 2 64 65 NOR
X69 en 63 66 NAND
X70 14 37 67 NOR
X71 48 67 68 NOR
X72 5 68 50.3 NOR
X73 34 39 69 NOR
X74 33 40 70 NAND
X75 cal_count.0 70 71 NAND
X76 cal_count.0 state.2 72 NAND
X77 47 72 73 NAND
X78 71 73 74.0 NAND
X79 cal_count.1 47 75 NOR
X80 cal_count.0 cal_count.1 76 NAND
X81 76 77 NOT
X82 comp 76 78 NAND
X83 comp 76 79 NOR
X84 6 77 80 NAND
X85 cal_count.0 cal_count.1 81 NOR
X86 78 80 82 NAND
X87 81 82 83 NOR
X88 comp 81 84 NAND
X89 69 84 85 NAND
X90 83 85 86 NOR
X91 75 86 74.1 NOR
X92 cal_count.2 47 87 NOR
X93 80 84 88 NAND
X94 7 88 89 NAND
X95 69 89 90 NAND
X96 7 88 91 NOR
X97 90 91 92 NOR
X98 87 92 74.2 NOR
X99 cal_count.3 48 93 NAND
X100 cal_count.2 79 94 NAND
X101 94 95 NOT
X102 cal_count.2 84 96 NOR
X103 96 97 NOT
X104 95 96 98 NOR
X105 94 97 99 NAND
X106 8 99 100 NAND
X107 cal_count.3 98 101 NAND
X108 100 101 102 NAND
X109 69 102 103 NAND
X110 93 103 74.3 NAND
X111 9 66 104 NAND
X112 33 42 105 NAND
X113 13 62 106 NOR
X114 state.1 61 107 NAND
X115 mask.0 107 108 NOR
X116 63 108 109 NOR
X117 105 109 110 NAND
X118 104 110 111 NAND
X119 9 31 112 NOR
X120 62 112 113 NAND
X121 111 113 114 NAND
X122 calibrate 29 115 NOR
X123 28 115 116 NOR
X124 34 40 117 NOR
X125 33 39 118 NAND
X126 trim_mask.0 117 119 NAND
X127 8 119 120 NOR
X128 trim_val.0 120 121 NOR
X129 116 121 122.0 NOR
X130 trim_mask.1 117 123 NAND
X131 8 123 124 NOR
X132 trim_val.1 124 125 NOR
X133 116 125 122.1 NOR
X134 trim_mask.2 117 126 NAND
X135 8 126 127 NOR
X136 trim_val.2 127 128 NOR
X137 116 128 122.2 NOR
X138 trim_mask.3 117 129 NAND
X139 8 129 130 NOR
X140 trim_val.3 130 131 NOR
X141 116 131 122.3 NOR
X142 trim_mask.4 117 132 NAND
X143 8 132 133 NOR
X144 14 25 134 NAND
X145 11 116 135 NOR
X146 133 135 136 NOR
X147 134 136 122.4 NAND
X148 calibrate 30 137 NAND
X149 34 137 138 NAND
X150 70 138 139 NAND
X151 trim_mask.0 139 140 NAND
X152 123 140 141.0 NAND
X153 trim_mask.1 139 142 NAND
X154 126 142 141.1 NAND
X155 trim_mask.2 139 143 NAND
X156 129 143 141.2 NAND
X157 trim_mask.3 139 144 NAND
X158 132 144 141.3 NAND
X159 trim_mask.4 118 145 NAND
X160 137 145 141.4 NAND
X161 mask.1 106 146 NAND
X162 31 45 147 NAND
X163 61 147 148 NAND
X164 mask.0 148 149 NAND
X165 146 149 150.0 NAND
X166 mask.2 106 151 NAND
X167 mask.1 148 152 NAND
X168 151 152 150.1 NAND
X169 mask.3 106 153 NAND
X170 mask.2 148 154 NAND
X171 153 154 150.2 NAND
X172 mask.4 106 155 NAND
X173 mask.3 148 156 NAND
X174 155 156 150.3 NAND
X175 mask.5 106 157 NAND
X176 mask.4 148 158 NAND
X177 157 158 150.4 NAND
*X178 mask.6 106 159 NAND
X179 mask.5 148 160 NAND
X180 106 160 150.5 NAND
*X181 mask.7 106 161 NAND
*X182 mask.6 148 162 NAND
*X183 161 162 150.6 NAND
*X184 mask.8 106 163 NAND
*X185 mask.7 148 164 NAND
*X186 163 164 150.7 NAND
*X187 mask.9 106 165 NAND
*X188 mask.8 148 166 NAND
*X189 165 166 150.8 NAND
*X190 mask.9 65 167 NOR
*X191 106 167 150.9 NOR
X192 25 27 168 NOR
X193 13 14 169 NOR
X194 state.1 state.2 170 NAND
X195 105 170 171 NAND
X196 state.0 171 172 NAND
X197 147 168 173 NAND
X198 108 173 174 NOR
X199 172 174 175.0 NAND
X200 65 108 176 NOR
X201 115 169 177 NOR
X202 176 177 175.1 NAND
X203 mask.0 106 178 NAND
X204 138 169 179 NOR
X205 178 179 175.2 NAND
X206 cal 65 180 NAND
X207 47 105 181 NAND
X208 calibrate 181 182 NAND
X209 180 182 183 NAND
X210 comp 106 184 NAND
X211 15 184 185 NAND
X212 mask.0 result.0 ctln.0 NOR
X213 ctln.0 ctlp.0 NOT
X214 185 ctlp.0 186 NAND
X215 65 186 187.0 NOR
X216 16 184 188 NAND
X217 mask.1 result.1 ctln.1 NOR
X218 ctln.1 ctlp.1 NOT
X219 188 ctlp.1 189 NAND
X220 65 189 187.1 NOR
X221 17 184 190 NAND
X222 mask.2 result.2 ctln.2 NOR
X223 ctln.2 ctlp.2 NOT
X224 190 ctlp.2 191 NAND
X225 65 191 187.2 NOR
X226 18 184 192 NAND
X227 mask.3 result.3 ctln.3 NOR
X228 ctln.3 ctlp.3 NOT
X229 192 ctlp.3 193 NAND
X230 65 193 187.3 NOR
X231 19 184 194 NAND
X232 mask.4 result.4 ctln.4 NOR
X233 ctln.4 ctlp.4 NOT
X234 194 ctlp.4 195 NAND
X235 65 195 187.4 NOR
X236 20 184 196 NAND
X237 mask.5 result.5 ctln.5 NOR
X238 ctln.5 ctlp.5 NOT
X239 196 ctlp.5 197 NAND
X240 65 197 187.5 NOR
*X241 21 184 198 NAND
*X242 mask.6 result.6 ctln.6 NOR
*X243 ctln.6 ctlp.6 NOT
*X244 198 ctlp.6 199 NAND
*X245 65 199 187.6 NOR
*X246 22 184 200 NAND
*X247 mask.7 result.7 ctln.7 NOR
*X248 ctln.7 ctlp.7 NOT
*X249 200 ctlp.7 201 NAND
*X250 65 201 187.7 NOR
*X251 23 184 202 NAND
*X252 mask.8 result.8 ctln.8 NOR
*X253 ctln.8 ctlp.8 NOT
*X254 202 ctlp.8 203 NAND
*X255 65 203 187.8 NOR
*X256 24 184 204 NAND
*X257 mask.9 result.9 ctln.9 NOR
*X258 ctln.9 ctlp.9 NOT
*X259 204 ctlp.9 205 NAND
*X260 65 205 187.9 NOR
X261 trim_mask.0 trim_val.0 trimb.0 NOR
X262 trimb.0 trim.0 NOT
X263 trim_val.1 trim_mask.1 trimb.1 NOR
X264 trimb.1 trim.1 NOT
X265 trim_val.2 trim_mask.2 trimb.2 NOR
X266 trimb.2 trim.2 NOT
X267 trim_val.3 trim_mask.3 trimb.3 NOR
X268 trimb.3 trim.3 NOT
X269 trim_val.4 trim_mask.4 trimb.4 NOR
X270 trimb.4 trim.4 NOT
X271 9 clk clkc NOR
X272 rstn 206 NOT
X273 rstn 207 NOT
X274 rstn 208 NOT
X275 rstn 209 NOT
X276 rstn 210 NOT
X277 rstn 211 NOT
X278 rstn 212 NOT
X279 rstn 213 NOT
X280 rstn 214 NOT
X281 rstn 215 NOT
X282 rstn 216 NOT
X283 rstn 217 NOT
X284 rstn 218 NOT
X285 rstn 219 NOT
X286 rstn 220 NOT
X287 rstn 221 NOT
X288 rstn 222 NOT
X289 rstn 223 NOT
X290 rstn 224 NOT
X291 rstn 225 NOT
X292 rstn 226 NOT
X293 rstn 227 NOT
X294 rstn 228 NOT
X295 rstn 229 NOT
X296 rstn 230 NOT
X297 rstn 231 NOT
X298 rstn 232 NOT
X299 rstn 233 NOT
X300 rstn 234 NOT
X301 rstn 235 NOT
X302 rstn 236 NOT
X303 rstn 237 NOT
X304 rstn 238 NOT
X305 rstn 239 NOT
X306 rstn 240 NOT
X307 rstn 241 NOT
X308 rstn 242 NOT
X309 rstn 243 NOT
X310 rstn 244 NOT
X311 rstn 245 NOT
X312 rstn 246 NOT
X313 rstn 247 NOT
X314 clk 187.0 result.0 0s 206 DFFSR
X315 clk 187.1 result.1 0s 207 DFFSR
X316 clk 187.2 result.2 0s 208 DFFSR
X317 clk 187.3 result.3 0s 209 DFFSR
X318 clk 187.4 result.4 0s 210 DFFSR
X319 clk 187.5 result.5 0s 211 DFFSR
*X320 clk 187.6 result.6 0s 212 DFFSR
*X321 clk 187.7 result.7 0s 213 DFFSR
*X322 clk 187.8 result.8 0s 214 DFFSR
*X323 clk 187.9 result.9 0s 215 DFFSR
X324 clk 183 calibrate 0s 216 DFFSR
X325 clk 175.0 state.0 0s 217 DFFSR
X326 clk 175.1 state.1 0s 218 DFFSR
X327 clk 175.2 state.2 0s 219 DFFSR
X328 clk 150.0 mask.0 0s 220 DFFSR
X329 clk 150.1 mask.1 0s 221 DFFSR
X330 clk 150.2 mask.2 0s 222 DFFSR
X331 clk 150.3 mask.3 0s 223 DFFSR
X332 clk 150.4 mask.4 0s 224 DFFSR
X333 clk 150.5 mask.5 0s 225 DFFSR
X334 clk 150.6 mask.6 0s 226 DFFSR
X335 clk 150.7 mask.7 0s 227 DFFSR
X336 clk 150.8 mask.8 0s 228 DFFSR
X337 clk 150.9 mask.9 0s 229 DFFSR
X338 clk 141.0 trim_mask.0 0s 230 DFFSR
X339 clk 141.1 trim_mask.1 0s 231 DFFSR
X340 clk 141.2 trim_mask.2 0s 232 DFFSR
X341 clk 141.3 trim_mask.3 0s 233 DFFSR
X342 clk 141.4 trim_mask.4 0s 234 DFFSR
X343 clk 122.0 trim_val.0 0s 235 DFFSR
X344 clk 122.1 trim_val.1 0s 236 DFFSR
X345 clk 122.2 trim_val.2 0s 237 DFFSR
X346 clk 122.3 trim_val.3 0s 238 DFFSR
X347 clk 122.4 trim_val.4 0s 239 DFFSR
X348 clk 114 en_co_clk 0s 240 DFFSR
X349 clk 74.0 cal_count.0 241 0s DFFSR
X350 clk 74.1 cal_count.1 242 0s DFFSR
X351 clk 74.2 cal_count.2 243 0s DFFSR
X352 clk 74.3 cal_count.3 0s 244 DFFSR
X353 clk 50.0 cal_itt.0 0s 245 DFFSR
X354 clk 50.1 cal_itt.1 0s 246 DFFSR
X355 clk 50.2 cal_itt.2 0s 247 DFFSR
X356 clk 50.3 cal_itt.3 0s 1 DFFSR
.ends sarlogic
